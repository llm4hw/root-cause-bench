----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11.03.2024 02:00:57
-- Design Name: 
-- Module Name: SignalVariableError - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top6 is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           out1 : out STD_LOGIC);
end top6;

architecture Behavioral of top6 is
    signal signal1 : STD_LOGIC := '0';
    variable variable1 : STD_LOGIC := '0';
begin
    process (clk, rst)
    begin
        if rst = '1' then
            signal1 <= '0';
            variable1 := '0'; 
        elsif rising_edge(clk) then
            variable1 := signal1;
        end if;
    end process;


    out1 <= signal1;
end Behavioral;

